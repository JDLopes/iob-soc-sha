`define OPCODE_W 2


